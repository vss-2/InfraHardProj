//Modulo simples o qual recebe como entrada 2 valores e sua saida e o XOR deles
module XORR (input logic sinal_1, sinal_2, output logic Xor_out);	
		assign Xor_out = sinal_1 ^ sinal_2;	
endmodule: XORR
